comparator_inst : comparator PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		ageb	 => ageb_sig
	);
