lpm_add_sub0_inst : lpm_add_sub0 PORT MAP (
		add_sub	 => add_sub_sig,
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		cout	 => cout_sig,
		result	 => result_sig
	);
