library IEEE; use IEEE.STD_LOGIC_1164.all;

entity mux4_12 is
  port (
    d0, d1, d2, d3 : in STD_LOGIC_VECTOR(11 downto 0);
    s : in STD_LOGIC_VECTOR(1 downto 0);
    y : out STD_LOGIC_VECTOR(11 downto 0)
  );
end mux4_12;

architecture synth of mux4_12 is
  component mux2
    generic (width : integer := 8);  --default value, if not given in "init"
    port (
      d0, d1 : in STD_LOGIC_VECTOR(width-1 downto 0);
      s : in STD_LOGIC;
      y : out STD_LOGIC_VECTOR(width-1 downto 0)
    );
  end component;

  signal lowb, highb: STD_LOGIC_VECTOR(11 downto 0);

begin
  -- for 4-8 mux
 -- lowmux: mux2 port map(d0, d1, s(0), low);
 -- highmux: mux2 port map(d2, d3, s(0), high);
  --outmux: mux2 port map(low, high, s(1), y);
  -- for 4-12 mux
  lowmux:   mux2 generic map(12)
                 port map(d0, d1, s(0), lowb);
  highmux:  mux2 generic map(12)
                 port map(d2, d3, s(0), highb);
  outmux:   mux2 generic map(12)
                 port map(lowb, highb, s(1), y);  
end synth; 