altfp_mult0_inst : altfp_mult0 PORT MAP (
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		overflow	 => overflow_sig,
		result	 => result_sig
	);
