library IEEE; use IEEE.STD_LOGIC_1164.all;

entity flopenr is
  port (
    clk, reset, en : in STD_LOGIC;
    d : in STD_LOGIC_VECTOR(3 downto 0);
    q : out STD_LOGIC_VECTOR(3 downto 0)
  );
end flopenr;

architecture synth of flopenr is
begin
  process (clk, reset, en) begin
    if reset then
      q <= "0000"; --similar to q <= (others => '0');
    elsif rising_edge(clk) then
      if en then
        q <= d;
      end if;  
    end if;
  end process;
end synth; 