-- Copyright (C) 1991-2011 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II"
-- VERSION		"Version 11.0 Build 208 07/03/2011 Service Pack 1 SJ Web Edition"
-- CREATED		"Sun Feb 14 17:11:50 2021"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY decoder_hex_7 IS 
	PORT
	(
		X0 :  IN  STD_LOGIC;
		X1 :  IN  STD_LOGIC;
		X2 :  IN  STD_LOGIC;
		X3 :  IN  STD_LOGIC;
		a :  OUT  STD_LOGIC;
		b :  OUT  STD_LOGIC;
		c :  OUT  STD_LOGIC;
		d :  OUT  STD_LOGIC;
		e :  OUT  STD_LOGIC;
		f :  OUT  STD_LOGIC;
		g :  OUT  STD_LOGIC
	);
END decoder_hex_7;

ARCHITECTURE bdf_type OF decoder_hex_7 IS 

SIGNAL	not_x0 :  STD_LOGIC;
SIGNAL	not_x0_nor_not_x1 :  STD_LOGIC;
SIGNAL	not_x1 :  STD_LOGIC;
SIGNAL	not_x1_nor_not_x2 :  STD_LOGIC;
SIGNAL	not_x2 :  STD_LOGIC;
SIGNAL	not_x2_nor_x3 :  STD_LOGIC;
SIGNAL	not_x3 :  STD_LOGIC;
SIGNAL	x1_nor_not_x2 :  STD_LOGIC;
SIGNAL	x1_nor_x2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;


BEGIN 



SYNTHESIZED_WIRE_0 <= NOT(not_x2_nor_x3 OR X0);


SYNTHESIZED_WIRE_18 <= NOT(SYNTHESIZED_WIRE_0 OR SYNTHESIZED_WIRE_1 OR not_x1_nor_not_x2 OR SYNTHESIZED_WIRE_2);


SYNTHESIZED_WIRE_8 <= NOT(not_x0_nor_not_x1 OR SYNTHESIZED_WIRE_3);


SYNTHESIZED_WIRE_34 <= NOT(not_x3 OR not_x0);


SYNTHESIZED_WIRE_3 <= NOT(X0 OR X1);


not_x0_nor_not_x1 <= NOT(not_x0 OR not_x1);


SYNTHESIZED_WIRE_37 <= NOT(not_x3 OR X1 OR not_x0);


c <= NOT(SYNTHESIZED_WIRE_4);



SYNTHESIZED_WIRE_4 <= NOT(SYNTHESIZED_WIRE_5 OR not_x2_nor_x3 OR SYNTHESIZED_WIRE_6);


SYNTHESIZED_WIRE_5 <= NOT(SYNTHESIZED_WIRE_7 OR X2);


SYNTHESIZED_WIRE_7 <= NOT(X3 OR not_x1);


SYNTHESIZED_WIRE_36 <= NOT(SYNTHESIZED_WIRE_8 OR X3);


SYNTHESIZED_WIRE_1 <= NOT(X1 OR X2 OR not_x3);


SYNTHESIZED_WIRE_6 <= NOT(not_x1_nor_not_x2 OR not_x0);


d <= NOT(SYNTHESIZED_WIRE_9);



SYNTHESIZED_WIRE_9 <= NOT(SYNTHESIZED_WIRE_10 OR SYNTHESIZED_WIRE_11 OR SYNTHESIZED_WIRE_12);


SYNTHESIZED_WIRE_11 <= NOT(SYNTHESIZED_WIRE_13 OR not_x2);


SYNTHESIZED_WIRE_13 <= NOT(SYNTHESIZED_WIRE_14 OR SYNTHESIZED_WIRE_15);


SYNTHESIZED_WIRE_12 <= NOT(not_x3 OR X1);


SYNTHESIZED_WIRE_14 <= NOT(not_x0 OR X1);


SYNTHESIZED_WIRE_15 <= NOT(not_x1 OR X0);


SYNTHESIZED_WIRE_10 <= NOT(X2 OR SYNTHESIZED_WIRE_16);


SYNTHESIZED_WIRE_16 <= NOT(not_x0_nor_not_x1 OR SYNTHESIZED_WIRE_17);


a <= NOT(SYNTHESIZED_WIRE_18);



SYNTHESIZED_WIRE_17 <= NOT(X0 OR X3);


SYNTHESIZED_WIRE_21 <= NOT(SYNTHESIZED_WIRE_19 OR SYNTHESIZED_WIRE_20);


SYNTHESIZED_WIRE_20 <= NOT(x1_nor_not_x2 OR X0);


x1_nor_not_x2 <= NOT(X1 OR not_x2);


SYNTHESIZED_WIRE_19 <= NOT(x1_nor_x2 OR not_x3);


e <= NOT(SYNTHESIZED_WIRE_21);



f <= NOT(SYNTHESIZED_WIRE_22);



g <= NOT(SYNTHESIZED_WIRE_23);



SYNTHESIZED_WIRE_22 <= NOT(SYNTHESIZED_WIRE_24 OR SYNTHESIZED_WIRE_25 OR SYNTHESIZED_WIRE_38);


not_x2_nor_x3 <= NOT(X3 OR not_x2);


SYNTHESIZED_WIRE_38 <= NOT(X3 OR not_x2 OR X1);


SYNTHESIZED_WIRE_30 <= NOT(X2 OR not_x1);


SYNTHESIZED_WIRE_25 <= NOT(x1_nor_not_x2 OR not_x3);


SYNTHESIZED_WIRE_23 <= NOT(SYNTHESIZED_WIRE_38 OR SYNTHESIZED_WIRE_28 OR SYNTHESIZED_WIRE_29);


SYNTHESIZED_WIRE_24 <= NOT(SYNTHESIZED_WIRE_30 OR X0);


SYNTHESIZED_WIRE_28 <= NOT(SYNTHESIZED_WIRE_31 OR not_x1);


SYNTHESIZED_WIRE_32 <= NOT(not_x2 OR X0);


SYNTHESIZED_WIRE_29 <= NOT(SYNTHESIZED_WIRE_32 OR not_x3);


SYNTHESIZED_WIRE_31 <= NOT(not_x2 OR not_x0);


not_x1 <= NOT(X1);



b <= NOT(SYNTHESIZED_WIRE_33);



not_x0 <= NOT(X0);



not_x1_nor_not_x2 <= NOT(not_x2 OR not_x1);


not_x2 <= NOT(X2);



SYNTHESIZED_WIRE_35 <= NOT(SYNTHESIZED_WIRE_34 OR X2);


not_x3 <= NOT(X3);



SYNTHESIZED_WIRE_2 <= NOT(not_x0 OR X3 OR x1_nor_x2);


x1_nor_x2 <= NOT(X2 OR X1);


SYNTHESIZED_WIRE_33 <= NOT(SYNTHESIZED_WIRE_35 OR SYNTHESIZED_WIRE_36 OR SYNTHESIZED_WIRE_37);


END bdf_type;